module decoder_4to16

	# (parameter N = 4)
	
	(input [N-1:0] 		   a,
	 output wire [2**N-1:0] d
	);
	
	decoder_3to8 DEC1 (
	.a(a[N-2:0]),
	.a3(~a[N-1]),
	.d(d[2**(N-1)-1:0])
	);

	decoder_3to8 DEC2 (
	.a(a[N-2:0]),
	.a3(a[N-1]),
	.d(d[2**N-1:2**(N-1)])
	);
	
endmodule